// Assignment 1
module Assignment_1();
  
  // Displays the message in the console on a new line with a TAB before
  initial begin
    $display("\n\t My Name is Praba and I start the course today jun 11th 2025 \n"); 
  end
  
endmodule